library verilog;
use verilog.vl_types.all;
entity tb_FinalCPU is
end tb_FinalCPU;
